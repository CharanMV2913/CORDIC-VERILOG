module Cordic (
    input clk,
    input ena,
    input [WIDTH-1:0] Xi,
    input [WIDTH-1:0] Yi,
    output reg [WIDTH + EXTEND_PRECISION -1:0] R,
    output reg [AWIDTH -1:0] A
);

parameter PIPELINE = 15;
parameter WIDTH = 16;
parameter AWIDTH = 16;
parameter EXTEND_PRECISION = 4;
parameter ANG = 20;
parameter PRECISION = WIDTH + EXTEND_PRECISION;

// Define types for arrays
typedef logic [PRECISION:0] XYVector [0:PIPELINE];
typedef logic [ANG-1:0] ZVector [0:PIPELINE];

// Define signals
reg [PRECISION:0] X [0:PIPELINE];
reg [PRECISION:0] Y [0:PIPELINE];
reg [ANG-1:0] Z [0:PIPELINE];

// Architecture body
initial begin
    // Fill first nodes
    X[0][PRECISION:EXTEND_PRECISION] = {1'b0, Xi}; // fill msb of X0
    for (int n = EXTEND_PRECISION - 1; n >= 0; n = n - 1) begin
        X[0][n] = 1'b0; // fill lsb with '0'
    end

    Y[0][PRECISION:EXTEND_PRECISION] = {Yi[WIDTH - 1], Yi}; // fill msb of Y0
    for (int n = EXTEND_PRECISION - 1; n >= 0; n = n - 1) begin
        Y[0][n] = 1'b0; // fill lsb with '0'
    end

    for (int n = ANG - 1; n >= 0; n = n - 1) begin
        Z[0][n] = 1'b0; // fill Z with '0'
    end

    // Generate pipeline
    for (int n = 1; n <= PIPELINE; n = n + 1) begin
        CordicPipe Pipe (
            .clk(clk),
            .ena(ena),
            .Xi(X[n-1]),
            .Yi(Y[n-1]),
            .Zi(Z[n-1]),
            .Xo(X[n]),
            .Yo(Y[n]),
            .Zo(Z[n])
        );
    end

    // Assign outputs
    R = X[PIPELINE][PRECISION-1:0];
    A = Z[PIPELINE][ANG-1:ANG-AWIDTH];
end

endmodule
